`ifndef _constants_sv_
`define _constants_sv_
/*
`define WORD_SIZE 32
`define TYPE_WIDTH 5
`define VALUE_WIDTH 13
define MEM_BYTES 8192
`define MEM_TOTAL `MEM_BYTES * `WORD_SIZE

// File I/O
`define EOF -1
`define ERR -2

`define MEM_ERR 32'bz

// Memory type *probably temporary until RAM gets used.*
typedef integer   addr_t;
*/
// Various types
//`define type_t [`TYPE_WIDTH:0]
//`define addr_t [`VALUE_WIDTH:0]
//`define bus_t [`WORD_SIZE:0]

`endif
