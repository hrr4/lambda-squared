module Computer(
		input  KEY[0], 
		output LEDR[0]
		);
   
   
   
   
endmodule
